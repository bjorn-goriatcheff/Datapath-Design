`include "CPU.v"

module CPU_fixture;
endmodule
