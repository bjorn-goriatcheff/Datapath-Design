module Registers(
	output reg[15:0] Data1,
	output reg[15:0] Data2,
	output reg[15:0] Data15,
	input [3:0] ReadAdd1,
	input [3:0] ReadAdd2,
	input [3:0] WriteReg1,
	input [3:0] WriteReg2,
	input WriteDst
);






endmodule
