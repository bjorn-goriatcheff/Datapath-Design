`include "PC.v"
`include "Adder2.v"
`include "INS.v"
`include "Registers.v"
`include "ALU.v"
`include "Sign.v"
`include "SignBr.v"
`include "Zero.v"
`include "MU3x1.v"
`include "MU4x1.v"
`include "ALU_CONTROL.v"
`include "CONTROL.v"
`include "Memory.v"
`include "AdderBr.v"
`include "SSL.v"
`include "XOR.v"
`include "CMP.v"
`include "BufferIFID.v"
`include "BufferIDEX.v"
`include "BufferEXMEM.v"
`include "BufferMEMWB.v"
`include "Forward.v"
`include "Gather.v"


module CPU;




endmodule
