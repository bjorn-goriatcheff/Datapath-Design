module CPU;
endmodule
